// Interface

// jkff_if.sv
interface jkff_if (input logic clk);
    logic rstn;
    logic j;
    logic k;
    logic q;
endinterface

