interface comp_if;
    logic [3:0] A;
    logic [3:0] B;
    logic A_gt_B;
    logic A_lt_B;
    logic A_eq_B;
endinterface

