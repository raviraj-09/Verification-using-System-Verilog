// Interface

interface srff_if (input logic clk);
    logic rstn;
    logic s;
    logic r;
    logic q;
endinterface

