
interface full_adder_if;
    logic a, b, cin;
    logic sum, carry;
endinterface
