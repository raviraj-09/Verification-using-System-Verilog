
interface half_adder_if;
    logic a, b;
    logic sum, carry;
endinterface
